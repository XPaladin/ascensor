program automatic test(algoritmo_io.TB algoritmo);
	initial begin
		$vcdpluson;
		reset();
	end
	task reset();
		# TODO!!!!!!!!!!!
	endtask
endprogram
