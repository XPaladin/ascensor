module ALGORITMO (solicitudes, cambio_piso, trabajando, estado_pisos, estado_ascensor, motor)
endmodule